domain KWGR614 broadcast
